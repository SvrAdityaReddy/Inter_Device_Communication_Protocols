module uartTest;
    
endmodule