module uart (
    
);
    
endmodule