module spi_master ();
    
endmodule

module spi_slave ();
    
endmodule
